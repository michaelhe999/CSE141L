module instruction_memory(
    input logic [31:0] pc,
    output logic [8:0] instruction
);

    always_comb begin
        instruction = //value at pc
    end
);

endmodule